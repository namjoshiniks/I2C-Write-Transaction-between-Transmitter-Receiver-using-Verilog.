module MockReciver(SDA);

inout SDA;
reg direction;
reg SDAAck;

//assign SDA = (direction) ? SDAAck : 1'bz;

endmodule

