module ShiftBuf1Reg_tb();

reg clk,signalShift,signalLoad;
reg [31:0] TxIn;
wire dout;
ShiftBuf1Reg MUT(clk,signalShift,signalLoad,TxIn,dout);

always
#5 clk = ~clk;

initial begin
clk = 1'b0;
signalShift = 1'b0;
signalLoad  = 1'b1;
TxIn = 14;

/*@(posedge clk)
begin
signalLoad = 1'b1;
end
*/
@(posedge clk)
begin
signalLoad = 1'b0;
signalShift = 1'b1;
end

@(posedge clk)
begin
signalLoad = 1'b0;
signalShift = 1'b1;
end

@(posedge clk)
begin
signalLoad = 1'b0;
signalShift = 1'b1;
end

@(posedge clk)
begin
signalLoad = 1'b0;
signalShift = 1'b1;
end

end
endmodule

